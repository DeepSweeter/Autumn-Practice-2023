interface interface_Intern (
    input Clk
);
    logic SampleData, TransferData;
endinterface